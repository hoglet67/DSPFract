library ieee;
use ieee.std_logic_1164.all;

package dsp_fractal_defs is

    subtype iterations_type is std_logic_vector(11 downto 0);

end package dsp_fractal_defs;
